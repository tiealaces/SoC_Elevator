
`define CLK_FREQ 100_000_000